module char_decoder(
		output reg [127:0] OUT,
		input [6:0] IN
	);
	always @(*)
	begin
		begin case(IN)
            7'd32: OUT = {128{1'b0}}; // space
            
            7'd48: OUT = {64'b00000000_00111000_01000100_01001100_01010100_
                            01010100_01100100_01000100_00111000, 56{1'b0}}; // '0'
            7'd49: OUT = {64'b00000000_00010000_00110000_01010000_00010000_
                            00010000_00010000_00010000_01111100, 56{1'b0}}; // '1'
            7'd50: OUT = {64'b00000000_00111000_01000100_00000100_00001000_
                            00010000_00100000_01000000_01111100, 56{1'b0}}; // '2'
            7'd51: OUT = {64'b00000000_00111000_01000100_00000100_00011000_
                            00000100_00000100_01000100_00111000, 56{1'b0}}; // '3'
            7'd52: OUT = {64'b00000000_00000100_00001100_00010100_00100100_
                            01000100_01111110_00000100_00000100, 56{1'b0}}; // '4'
            7'd53: OUT = {64'b00000000_01111100_01000000_01000000_01111000_
                            00000100_00000100_01000100_00111000, 56{1'b0}}; // '5'
            7'd54: OUT = {64'b00000000_00011000_00100000_01000000_01111000_
                            01000100_01000100_01000100_00111000, 56{1'b0}}; // '6'
            7'd55: OUT = {64'b00000000_01111100_00000100_00001000_00001000_
                            00010000_00010000_00100000_00100000, 56{1'b0}}; // '7'
            7'd56: OUT = {64'b00000000_00111000_01000100_01000100_00111000_
                            01000100_01000100_01000100_00111000, 56{1'b0}}; // '8'
            7'd56: OUT = {64'b00000000_00111000_01000100_01000100_01000100_
                            00111100_00000100_00001000_00110000, 56{1'b0}}; // '9'

			7'd65: OUT = {64'b00000000_00011000_00011000_00100100_00100100_
                            00111100_01000010_01000010_01000010, 56{1'b0}}; // 'A'
            7'd66: OUT = {64'b00000000_01111000_01000100_01000100_01111100_
                            01000010_01000010_01000010_01111100, 56{1'b0}}; // 'B'
			7'd67: OUT = {64'b00000000_00011100_00100010_01000000_01000000_
                            01000000_01000000_00100010_00011100, 56{1'b0}}; // 'C'
			7'd68: OUT = {64'b00000000_01111000_01000100_01000010_01000010_
                            01000010_01000010_01000100_01111000, 56{1'b0}}; // 'D'
			7'd69: OUT = {64'b00000000_01111110_01000000_01000000_01111000_
                            01000000_01000000_01000000_01111110, 56{1'b0}}; // 'E'
			7'd70: OUT = {64'b00000000_01111110_01000000_01000000_01111000_
                            01000000_01000000_01000000_01000000, 56{1'b0}}; // 'F'
			7'd71: OUT = {64'b00000000_00011100_00100010_01000000_01000000_
                            01001110_01000010_00100010_00011100, 56{1'b0}}; // 'G'
			7'd72: OUT = {64'b00000000_01000010_01000010_01000010_01111110_
                            01000010_01000010_01000010_01000010, 56{1'b0}}; // 'H'
			7'd73: OUT = {64'b00000000_00111000_00010000_00010000_00010000_
                            00010000_00010000_00010000_00111000, 56{1'b0}}; // 'I'
			7'd74: OUT = {64'b00000000_00001110_00000010_00000010_00000010_
                            00000010_00000010_00000010_00011110, 56{1'b0}}; // 'J'
			7'd75: OUT = {64'b00000000_01000010_01000100_01001000_01010000_
                            01110000_01001000_01000100_01000010, 56{1'b0}}; // 'K'
			7'd76: OUT = {64'b00000000_01000000_01000000_01000000_01000000_
                            01000000_01000000_01000000_01111110, 56{1'b0}}; // 'L'
			7'd77: OUT = {64'b00000000_11000110_11000110_10101010_10101010_
                            10010010_10010010_10000010_10000010, 56{1'b0}}; // 'M'
			7'd78: OUT = {64'b00000000_01100010_01100010_01010010_01010010_
                            01001010_01001010_01000110_01000110, 56{1'b0}}; // 'N'
			7'd79: OUT = {64'b00000000_00011000_00100100_01000100_01000100_
                            01000100_01000100_00100100_00011000, 56{1'b0}}; // 'O'
			7'd80: OUT = {64'b00000000_01111000_01000100_01000100_01000100_
                            01111000_01000000_01000000_01000000, 56{1'b0}}; // 'P'
			7'd81: OUT = {64'b00000000_00011000_00100100_01000100_01000100_
                            01000100_01000100_00100100_00011010_00000010, 48{1'b0}}; // 'Q'
			7'd82: OUT = {64'b00000000_01111000_01000100_01000100_01000100_
                            01111000_01001000_01000100_01000010, 56{1'b0}}; // 'R'
			7'd83: OUT = {64'b00000000_00111100_01000010_01000000_00110000_
                            00001100_00000010_01000010_00111100, 56{1'b0}}; // 'S'
			7'd84: OUT = {64'b00000000_11111110_00010000_00010000_00010000_
                            00010000_00010000_00010000_00010000, 56{1'b0}}; // 'T'
			7'd85: OUT = {64'b00000000_01000010_01000010_01000010_01000010_
                            01000010_01000010_01000010_00111100, 56{1'b0}}; // 'U'
			7'd86: OUT = {64'b00000000_10000010_10000010_01000100_01000100_
                            00101000_00101000_00010000_00010000, 56{1'b0}}; // 'V'
			7'd87: OUT = {64'b00000000_10000010_10010010_10010010_10101010_
                            10101010_01101100_01000100_01000100, 56{1'b0}}; // 'W'
			7'd88: OUT = {64'b00000000_01000010_01000010_00100100_00011000_
                            00011000_00100100_01000010_01000010, 56{1'b0}}; // 'Y'
            7'd89: OUT = {64'b00000000_10000010_10000010_01000100_00101000_
                            00010000_00010000_00010000_00010000, 56{1'b0}}; // 'X'
            7'd90: OUT = {64'b00000000_01111110_00000010_00000100_00001000_
                            00010000_00100000_01000000_01111110, 56{1'b0}}; // 'Z'
		endcase
	end
end module