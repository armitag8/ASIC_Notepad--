module char_decoder(
        output reg [127:0] OUT,
        input [6:0] IN
    );
    always @(*)
    begin
        case(IN[6:0])
            7'd32: OUT = {128{1'b0}}; // space
            7'd33: OUT = { {8{1'b0}}, {6{8'b00010000}}, 8'b00000000, 8'b00010000, {56{1'b0}}}; // "!"
            7'd34: OUT = {24'b00010100_00010100_00101000, {104{1'b0}}}; // '"'
            7'd35: OUT = {72'b00000000_00010100_00010100_01111110_00101000_00101000_11111100_01010000_01010000, {56{1'b0}}}; // "#"
            7'd36: OUT = {72'b00000000_00010000_00111100_01010000_01010000_00111000_00010100_00010100_01111000_00010000, {56{1'b0}}}; // "$"
            7'd37: OUT = {72'b00000000_01000100_10101000_10101000_01010000_00010100_00101010_00101010_01000100, {56{1'b0}}}; // "%"
            7'd38: OUT = {72'b00000000_00110000_01001000_01001000_00110010_01001010_01000100_01000100_00111010, {56{1'b0}}}; // "&"
            7'd39: OUT = {24'b00001000_00001000_00010000, {104{1'b0}}};// "'" single quote
            7'd40: OUT = {88'b00001000_00010000_00010000_00100000_00100000_00100000_00100000_00100000_00010000_00010000_00001000, {40{1'b0}}}; // "("
            7'd41: OUT = {88'b00100000_00010000_00010000_00001000_00001000_00001000_00001000_00001000_00010000_00010000_00100000, {40{1'b0}}}; // ")"
            7'd42: OUT = {{24{1'b0}}, 40'b00010000_01010100_00111000_01010100_00010000, {64{1'b0}}}; // "*" 
            7'd43: OUT = {{16{1'b0}}, 40'b00010000_00010000_01111100_00010000_00010000, {72{1'b0}}}; // "+"
            7'd44: OUT = {{56{1'b0}}, 32'b00001000_00001000_00001000_00010000,{40{1'b0}}}; // ','
            7'd45: OUT = {{40{1'b0}}, 8'b00111100 , {80{1'b0}}};// '-'
            7'd46: OUT = {{56{1'b0}}, 16'b00010000_00010000, {56{1'b0}}};// '.'
            7'd47: OUT = {80'b00000100_00000100_00001000_00001000_00010000_00010000_00100000_00100000_01000000_01000000, {48{1'b0}}};// '/'
            7'd48: OUT = {72'b00000000_00111000_01000100_01001100_01010100_01010100_01100100_01000100_00111000, {56{1'b0}}}; // '0'
            7'd49: OUT = {72'b00000000_00010000_00110000_01010000_00010000_00010000_00010000_00010000_01111100, {56{1'b0}}}; // '1'
            7'd50: OUT = {72'b00000000_00111000_01000100_00000100_00001000_00010000_00100000_01000000_01111100, {56{1'b0}}}; // '2'
            7'd51: OUT = {72'b00000000_00111000_01000100_00000100_00011000_00000100_00000100_01000100_00111000, {56{1'b0}}}; // '3'
            7'd52: OUT = {72'b00000000_00000100_00001100_00010100_00100100_01000100_01111110_00000100_00000100, {56{1'b0}}}; // '4'
            7'd53: OUT = {72'b00000000_01111100_01000000_01000000_01111000_00000100_00000100_01000100_00111000, {56{1'b0}}}; // '5'
            7'd54: OUT = {72'b00000000_00011000_00100000_01000000_01111000_01000100_01000100_01000100_00111000, {56{1'b0}}}; // '6'
            7'd55: OUT = {72'b00000000_01111100_00000100_00001000_00001000_00010000_00010000_00100000_00100000, {56{1'b0}}}; // '7'
            7'd56: OUT = {72'b00000000_00111000_01000100_01000100_00111000_01000100_01000100_01000100_00111000, {56{1'b0}}}; // '8'
            7'd57: OUT = {72'b00000000_00111000_01000100_01000100_01000100_00111100_00000100_00001000_00110000, {56{1'b0}}}; // '9'
            7'd58: OUT = {{24{1'b0}}, 40'b00010000_00010000_00000000_00010000_00010000, {64{1'b0}}}; // ":"
            7'd59: OUT = {88'b00000000_00000000_00000000_00001000_00001000_00000000_00000000_00001000_00001000_00001000_00010000, {40{1'b0}}};// ';'
            7'd60: OUT = {{24{1'b0}}, 40'b00000110_00011000_01100000_00011000_00000110, {64{1'b0}}}; // "<"
            7'd61: OUT = {{32{1'b0}}, 24'b01111110_00000000_01111110, {72{1'b0}}};// '='
            7'd62: OUT = {{24{1'b0}}, 40'b01100000_00011000_00000110_00011000_01100000, {64{1'b0}}}; // ">"
            7'd63: OUT = {72'b00000000_00111000_01000100_00000100_00001000_00010000_0001000_00000000_00001000, {56{1'b0}}}; // "?"
            7'd64: OUT = {{8{1'b0}}, 64'b00111000_01000100_10011010_10101010_10101010_10011100_01000000_00111101, {56{1'b0}}}; // "@"
            7'd65: OUT = {72'b00000000_00011000_00011000_00100100_00100100_00111100_01000010_01000010_01000010, {56{1'b0}}}; // 'A'
            7'd66: OUT = {72'b00000000_01111000_01000100_01000100_01111100_01000010_01000010_01000010_01111100, {56{1'b0}}}; // 'B'
            7'd67: OUT = {72'b00000000_00011100_00100010_01000000_01000000_01000000_01000000_00100010_00011100, {56{1'b0}}}; // 'C'
            7'd68: OUT = {72'b00000000_01111000_01000100_01000010_01000010_01000010_01000010_01000100_01111000, {56{1'b0}}}; // 'D'
            7'd69: OUT = {72'b00000000_01111110_01000000_01000000_01111000_01000000_01000000_01000000_01111110, {56{1'b0}}}; // 'E'
            7'd70: OUT = {72'b00000000_01111110_01000000_01000000_01111000_01000000_01000000_01000000_01000000, {56{1'b0}}}; // 'F'
            7'd71: OUT = {72'b00000000_00011100_00100010_01000000_01000000_01001110_01000010_00100010_00011100, {56{1'b0}}}; // 'G'
            7'd72: OUT = {72'b00000000_01000010_01000010_01000010_01111110_01000010_01000010_01000010_01000010, {56{1'b0}}}; // 'H'
            7'd73: OUT = {72'b00000000_00111000_00010000_00010000_00010000_00010000_00010000_00010000_00111000, {56{1'b0}}}; // 'I'
            7'd74: OUT = {72'b00000000_00001110_00000010_00000010_00000010_00000010_00000010_00000010_00011110, {56{1'b0}}}; // 'J'
            7'd75: OUT = {72'b00000000_01000010_01000100_01001000_01010000_01110000_01001000_01000100_01000010, {56{1'b0}}}; // 'K'
            7'd76: OUT = {72'b00000000_01000000_01000000_01000000_01000000_01000000_01000000_01000000_01111110, {56{1'b0}}}; // 'L'
            7'd77: OUT = {72'b00000000_11000110_11000110_10101010_10101010_10010010_10010010_10000010_10000010, {56{1'b0}}}; // 'M'
            7'd78: OUT = {72'b00000000_01100010_01100010_01010010_01010010_01001010_01001010_01000110_01000110, {56{1'b0}}}; // 'N'
            7'd79: OUT = {72'b00000000_00011000_00100100_01000010_01000010_01000010_01000010_00100100_00011000, {56{1'b0}}}; // 'O'
            7'd80: OUT = {72'b00000000_01111000_01000100_01000100_01000100_01111000_01000000_01000000_01000000, {56{1'b0}}}; // 'P'
            7'd81: OUT = {80'b00000000_00011000_00100100_01000010_01000010_01000010_01000010_00100100_00011010_00000010, {48{1'b0}}}; // 'Q'
            7'd82: OUT = {72'b00000000_01111000_01000100_01000100_01000100_01111000_01001000_01000100_01000010, {56{1'b0}}}; // 'R'
            7'd83: OUT = {72'b00000000_00111100_01000010_01000000_00110000_00001100_00000010_01000010_00111100, {56{1'b0}}}; // 'S'
            7'd84: OUT = {72'b00000000_11111110_00010000_00010000_00010000_00010000_00010000_00010000_00010000, {56{1'b0}}}; // 'T'
            7'd85: OUT = {72'b00000000_01000010_01000010_01000010_01000010_01000010_01000010_01000010_00111100, {56{1'b0}}}; // 'U'
            7'd86: OUT = {72'b00000000_10000010_10000010_01000100_01000100_00101000_00101000_00010000_00010000, {56{1'b0}}}; // 'V'
            7'd87: OUT = {72'b00000000_10000010_10010010_10010010_10101010_10101010_01101100_01000100_01000100, {56{1'b0}}}; // 'W'
            7'd88: OUT = {72'b00000000_01000010_01000010_00100100_00011000_00011000_00100100_01000010_01000010, {56{1'b0}}}; // 'X'
            7'd89: OUT = {72'b00000000_10000010_10000010_01000100_00101000_00010000_00010000_00010000_00010000, {56{1'b0}}}; // 'Y'
            7'd90: OUT = {72'b00000000_01111110_00000010_00000100_00001000_00010000_00100000_01000000_01111110, {56{1'b0}}}; // 'Z'
            7'd91: OUT = {88'b00111000_00100000_00100000_00100000_00100000_00100000_00100000_00100000_00100000_00100000_00111000, {40{1'b0}}};// '['
            7'd92: OUT = {80'b01000000_01000000_00100000_00100000_00010000_00010000_00001000_00001000_00000100_00000100, {48{1'b0}}};// '\'
            7'd93: OUT = {88'b00111000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00001000_00111000, {40{1'b0}}};// ']'
            7'd94: OUT = {48'b00010000_00010000_00101000_00101000_01000100_01000100, {80{1'b0}}}; // "^"
            7'd95: OUT = {{72{1'b0}}, 8'b11111110, {48{1'b0}}}; // "_"    
            7'd96: OUT =   {16'b00010000_00001000, {112{1'b0}}};// '`'  
            
            7'd97: OUT = {72'b00000000_00000000_00000000_00111000_00000100_00111100_01000100_01000100_00111100, {56{1'b0}}}; // 'a'
            7'd98: OUT = {72'b00000000_01000000_01000000_01111000_01000100_01000100_01000100_01000100_01111000, {56{1'b0}}}; // 'b'
            7'd99: OUT = {72'b00000000_00000000_00000000_00111000_01000100_01000000_01000000_01000100_00111000, {56{1'b0}}}; // 'c'
            7'd100: OUT = {72'b00000000_00000100_00000100_00111100_01000100_01000100_01000100_01000100_00111100, {56{1'b0}}}; // 'd'
            7'd101: OUT = {72'b00000000_00000000_00000000_00111000_01000100_01111100_01000000_01000100_00111000, {56{1'b0}}}; // 'e'
            7'd102: OUT = {72'b00000000_00011100_00100000_00100000_01111000_00100000_00100000_00100000_00100000, {56{1'b0}}}; // 'f'
            7'd103: OUT = {96'b00000000_00000000_00000000_00110100_01001000_01001000_00110000_01000000_00111100_01000010_01000010_00111100, {32{1'b0}}}; // 'g'
            7'd104: OUT = {72'b00000000_01000000_01000000_01000000_01110000_01001000_01001000_01001000_01001000, {56{1'b0}}}; // 'h'
            7'd105: OUT = {72'b00000000_00000000_00010000_00000000_00110000_00010000_00010000_00010000_00010000, {56{1'b0}}}; // 'i'
            7'd106: OUT = {88'b00000000_00000000_00000100_00000000_00001100_00000100_00000100_00000100_00000100_00000100_00111000, {40{1'b0}}}; // 'j'
            7'd107: OUT = {72'b00000000_01000000_01000000_01000100_01001000_01010000_01110000_01001000_01000100, {56{1'b0}}}; // 'k'
            7'd108: OUT = {72'b00000000_00110000_00010000_00010000_00010000_00010000_00010000_00010000_00001000, {56{1'b0}}}; // 'l'
            7'd109: OUT = {72'b00000000_00000000_00000000_01101000_01010100_01010100_01010100_01010100_01010100, {56{1'b0}}}; // 'm'
            7'd110: OUT = {72'b00000000_00000000_00000000_01111000_01000100_01000100_01000100_01000100_01000100, {56{1'b0}}}; // 'n'
            7'd111: OUT = {72'b00000000_00000000_00000000_00111000_01000100_01000100_01000100_01000100_00111000, {56{1'b0}}}; // 'O'
            7'd112: OUT = {96'b00000000_00000000_00000000_01111000_01000100_01000100_01000100_01000100_01111000_01000000_01000000_01000000, {32{1'b0}}}; // 'p'
            7'd113: OUT = {96'b00000000_00000000_00000000_00111100_01000100_01000100_01000100_01000100_00111100_00000100_00000100_00000100, {32{1'b0}}}; // 'q'
            7'd114: OUT = {72'b00000000_00000000_00000000_01011000_01100100_01000000_01000000_01000000_01000000, {56{1'b0}}}; // 'r'
            7'd115: OUT = {72'b00000000_00000000_00000000_00111100_01000000_00110000_00001000_00000100_01111000, {56{1'b0}}}; // 's'
            7'd116: OUT = {72'b00000000_01000000_01000000_01111000_01000000_01000000_01000000_01000000_00111000, {56{1'b0}}}; // 't'
            7'd117: OUT = {72'b00000000_00000000_00000000_01000100_01000100_01000100_01000100_01000100_00111100, {56{1'b0}}}; // 'u'
            7'd118: OUT = {72'b00000000_00000000_00000000_01000100_01000100_00101000_00101000_00010000_00010000, {56{1'b0}}}; // 'v'
            7'd119: OUT = {72'b00000000_00000000_00000000_01000100_01010100_01010100_01010100_00101000_00101000, {56{1'b0}}}; // 'w'
            7'd120: OUT = {72'b00000000_00000000_00000000_01000100_00101000_00010000_00010000_00101000_01000100, {56{1'b0}}}; // 'x'
            7'd121: OUT = {96'b00000000_00000000_00000000_01000100_01000100_00101000_00101000_00101000_00010000_00010000_00010000_00100000, {32{1'b0}}}; // 'y'
            7'd122: OUT = {72'b00000000_00000000_00000000_01111100_00000100_00001000_00010000_00100000_01111100, {56{1'b0}}}; // 'z'
            7'd123: OUT = {88'b00001100_00010000_00010000_00010000_00010000_01100000_00010000_00010000_00010000_00010000_00001100, {40{1'b0}}};// "{"
            7'd124: OUT = {{11{8'b00010000}}, {40{1'b0}}}; // "|"
            7'd125: OUT = {88'b01100000_00010000_00010000_00010000_00010000_00001100_00010000_00010000_00010000_00010000_01100000, {40{1'b0}}}; // "}"
            7'd126: OUT = {{32{1'b0}}, 16'b01110010_10011100, {80{1'b0}}}; // '~'
            
            default: OUT = {128{1'b0}}; // space AKA blank
        endcase
    end
endmodule
